library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity MUX_intf is
	port(
		  DATA_IN 		: IN STD_LOGIC_VECTOR(7 downto 0);
		  CONSTANT_BUS : IN STD_LOGIC_VECTOR(7 downto 0);
		  RAM_DATA_OUT_BUS: IN STD_LOGIC_VECTOR(7 downto 0);
		  IN_SEL				: IN STD_LOGIC_VECTOR(1 downto 0);
		  IN_SEL_OUT_BUS : OUT  std_logic_vector(7 downto 0)
		  );
end MUX_intf;

architecture MUX_arch of MUX_intf is

begin
INSEL_A_MUX : process(DATA_IN, CONSTANT_BUS, RAM_DATA_OUT_BUS, IN_SEL)
	 begin
		if(IN_SEL = "00") then
			IN_SEL_OUT_BUS <= DATA_IN;
		elsif(IN_SEL = "01") then
			IN_SEL_OUT_BUS <= RAM_DATA_OUT_BUS;
		else
			IN_SEL_OUT_BUS <= CONSTANT_BUS;
		end if;
	 end process INSEL_A_MUX;
end MUX_arch;